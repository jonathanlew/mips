`define opWidth 6
`define regWidth 5
`define immWidth 16
`define valWidth 32
`define PCWidth 9

//module decodeStage (//inputs
